-- GENERATED WITH MATLAB...

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package GOLAY_SEQ_pkg is 

	 constant GOLAY_A : std_logic_vector(0 to 128-1) := ( "01011001110000000101011011001111101001100011111101010110110011110101100111000000010101101100111101011001110000001010100100110000"); 
 
	 constant GOLAY_B : std_logic_vector(0 to 128-1) := ( "10100110001111111010100100110000010110011100000010101001001100000101100111000000010101101100111101011001110000001010100100110000"); 
 
end GOLAY_SEQ_pkg; 
